version 60
