hello

task phase2;
    display("phase2");
endtask
